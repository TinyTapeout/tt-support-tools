VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_logo_corner
  CLASS BLOCK ;
  FOREIGN tt_logo_corner ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  OBS
      LAYER TopMetal2 ;
        RECT 45.000 99.500 55.000 100.000 ;
        RECT 41.500 99.000 58.500 99.500 ;
        RECT 39.000 98.500 61.000 99.000 ;
        RECT 37.000 98.000 63.000 98.500 ;
        RECT 35.000 97.500 65.000 98.000 ;
        RECT 33.500 97.000 66.500 97.500 ;
        RECT 32.500 96.500 67.500 97.000 ;
        RECT 31.000 96.000 69.000 96.500 ;
        RECT 30.000 95.500 70.000 96.000 ;
        RECT 29.000 95.000 71.000 95.500 ;
        RECT 28.000 94.500 72.500 95.000 ;
        RECT 26.500 94.000 73.000 94.500 ;
        RECT 26.000 93.500 74.000 94.000 ;
        RECT 25.000 93.000 75.000 93.500 ;
        RECT 24.000 92.500 76.000 93.000 ;
        RECT 23.500 92.000 47.000 92.500 ;
        RECT 53.000 92.000 76.500 92.500 ;
        RECT 22.500 91.500 43.000 92.000 ;
        RECT 57.000 91.500 77.500 92.000 ;
        RECT 22.000 91.000 40.500 91.500 ;
        RECT 59.500 91.000 78.000 91.500 ;
        RECT 21.000 90.500 38.500 91.000 ;
        RECT 61.500 90.500 79.000 91.000 ;
        RECT 20.500 90.000 37.000 90.500 ;
        RECT 63.000 90.000 79.500 90.500 ;
        RECT 19.500 89.500 35.500 90.000 ;
        RECT 64.500 89.500 80.500 90.000 ;
        RECT 19.000 89.000 34.000 89.500 ;
        RECT 66.000 89.000 81.000 89.500 ;
        RECT 18.500 88.500 33.000 89.000 ;
        RECT 67.000 88.500 81.500 89.000 ;
        RECT 18.000 88.000 32.000 88.500 ;
        RECT 68.000 88.000 82.000 88.500 ;
        RECT 17.500 87.500 31.000 88.000 ;
        RECT 69.000 87.500 82.500 88.000 ;
        RECT 16.500 87.000 30.000 87.500 ;
        RECT 70.000 87.000 83.500 87.500 ;
        RECT 16.000 86.500 29.000 87.000 ;
        RECT 71.000 86.500 84.000 87.000 ;
        RECT 15.500 86.000 28.000 86.500 ;
        RECT 72.000 86.000 84.500 86.500 ;
        RECT 15.000 85.500 27.500 86.000 ;
        RECT 72.500 85.500 85.000 86.000 ;
        RECT 14.500 85.000 26.500 85.500 ;
        RECT 73.500 85.000 85.500 85.500 ;
        RECT 14.000 84.500 26.000 85.000 ;
        RECT 74.000 84.500 86.000 85.000 ;
        RECT 13.500 84.000 25.000 84.500 ;
        RECT 75.000 84.000 86.500 84.500 ;
        RECT 13.000 83.500 24.500 84.000 ;
        RECT 75.500 83.500 87.000 84.000 ;
        RECT 12.500 83.000 24.000 83.500 ;
        RECT 76.000 83.000 87.500 83.500 ;
        RECT 12.500 82.500 23.000 83.000 ;
        RECT 77.000 82.500 87.500 83.000 ;
        RECT 12.000 82.000 22.500 82.500 ;
        RECT 77.500 82.000 88.000 82.500 ;
        RECT 11.500 81.500 22.000 82.000 ;
        RECT 78.000 81.500 88.500 82.000 ;
        RECT 11.000 81.000 21.500 81.500 ;
        RECT 78.500 81.000 89.000 81.500 ;
        RECT 10.500 80.000 21.000 81.000 ;
        RECT 79.000 80.500 89.500 81.000 ;
        RECT 79.500 80.000 90.000 80.500 ;
        RECT 10.000 79.500 21.000 80.000 ;
        RECT 80.000 79.500 90.000 80.000 ;
        RECT 9.500 79.000 21.000 79.500 ;
        RECT 80.500 79.000 90.500 79.500 ;
        RECT 9.000 78.000 59.500 79.000 ;
        RECT 81.000 78.500 91.000 79.000 ;
        RECT 81.500 78.000 91.000 78.500 ;
        RECT 8.500 77.500 59.500 78.000 ;
        RECT 82.000 77.500 91.500 78.000 ;
        RECT 8.000 76.500 59.500 77.500 ;
        RECT 82.500 77.000 92.000 77.500 ;
        RECT 7.500 76.000 59.500 76.500 ;
        RECT 83.000 76.500 92.000 77.000 ;
        RECT 83.000 76.000 92.500 76.500 ;
        RECT 7.000 75.000 59.500 76.000 ;
        RECT 83.500 75.500 93.000 76.000 ;
        RECT 84.000 75.000 93.000 75.500 ;
        RECT 6.500 74.000 59.500 75.000 ;
        RECT 84.500 74.000 93.500 75.000 ;
        RECT 6.000 73.000 59.500 74.000 ;
        RECT 85.000 73.500 94.000 74.000 ;
        RECT 5.500 72.000 59.500 73.000 ;
        RECT 85.500 73.000 94.000 73.500 ;
        RECT 85.500 72.500 94.500 73.000 ;
        RECT 86.000 72.000 94.500 72.500 ;
        RECT 5.000 71.000 59.500 72.000 ;
        RECT 86.500 71.000 95.000 72.000 ;
        RECT 4.500 70.000 59.500 71.000 ;
        RECT 87.000 70.000 95.500 71.000 ;
        RECT 4.000 69.000 59.500 70.000 ;
        RECT 87.500 69.000 96.000 70.000 ;
        RECT 3.500 67.500 59.500 69.000 ;
        RECT 88.000 68.000 96.500 69.000 ;
        RECT 3.000 65.500 59.500 67.500 ;
        RECT 88.500 67.500 96.500 68.000 ;
        RECT 88.500 67.000 97.000 67.500 ;
        RECT 89.000 66.500 97.000 67.000 ;
        RECT 89.000 66.000 97.500 66.500 ;
        RECT 1.000 58.500 8.500 61.000 ;
        RECT 0.500 57.000 8.500 58.500 ;
        RECT 0.500 55.000 8.000 57.000 ;
        RECT 0.000 53.000 8.000 55.000 ;
        RECT 30.000 54.500 45.000 65.500 ;
        RECT 89.500 65.000 97.500 66.000 ;
        RECT 89.500 64.500 98.000 65.000 ;
        RECT 90.000 63.000 98.000 64.500 ;
        RECT 90.500 61.500 98.500 63.000 ;
        RECT 91.000 61.000 98.500 61.500 ;
        RECT 91.000 59.500 99.000 61.000 ;
        RECT 91.500 58.500 99.000 59.500 ;
        RECT 91.500 57.000 99.500 58.500 ;
        RECT 92.000 55.000 99.500 57.000 ;
        RECT 0.000 47.000 7.500 53.000 ;
        RECT 0.000 45.000 8.000 47.000 ;
        RECT 0.500 43.000 8.000 45.000 ;
        RECT 0.500 41.500 8.500 43.000 ;
        RECT 1.000 40.500 8.500 41.500 ;
        RECT 30.000 41.000 82.500 54.500 ;
        RECT 92.000 52.500 100.000 55.000 ;
        RECT 92.500 47.500 100.000 52.500 ;
        RECT 92.000 45.500 100.000 47.500 ;
        RECT 92.000 43.000 99.500 45.500 ;
        RECT 91.500 41.500 99.500 43.000 ;
        RECT 1.000 39.000 9.000 40.500 ;
        RECT 1.500 38.500 9.000 39.000 ;
        RECT 1.500 37.000 9.500 38.500 ;
        RECT 2.000 36.500 9.500 37.000 ;
        RECT 2.000 35.500 10.000 36.500 ;
        RECT 2.000 35.000 10.500 35.500 ;
        RECT 2.500 34.000 10.500 35.000 ;
        RECT 2.500 33.500 11.000 34.000 ;
        RECT 3.000 33.000 11.000 33.500 ;
        RECT 3.000 32.500 11.500 33.000 ;
        RECT 3.500 32.000 11.500 32.500 ;
        RECT 3.500 31.000 12.000 32.000 ;
        RECT 30.000 31.500 45.000 41.000 ;
        RECT 53.000 40.500 68.500 41.000 ;
        RECT 91.500 40.500 99.000 41.500 ;
        RECT 4.000 30.000 12.500 31.000 ;
        RECT 4.500 29.000 13.000 30.000 ;
        RECT 4.500 28.500 13.500 29.000 ;
        RECT 5.000 28.000 13.500 28.500 ;
        RECT 5.000 27.500 14.000 28.000 ;
        RECT 5.500 26.500 14.500 27.500 ;
        RECT 6.000 26.000 15.000 26.500 ;
        RECT 6.500 25.000 15.500 26.000 ;
        RECT 7.000 24.500 16.000 25.000 ;
        RECT 7.000 24.000 16.500 24.500 ;
        RECT 7.500 23.500 17.000 24.000 ;
        RECT 8.000 23.000 17.000 23.500 ;
        RECT 8.000 22.500 17.500 23.000 ;
        RECT 8.500 22.000 18.000 22.500 ;
        RECT 9.000 21.500 18.500 22.000 ;
        RECT 9.000 21.000 19.000 21.500 ;
        RECT 9.500 20.500 19.500 21.000 ;
        RECT 10.000 20.000 20.000 20.500 ;
        RECT 10.000 19.500 20.500 20.000 ;
        RECT 10.500 19.000 21.000 19.500 ;
        RECT 11.000 18.500 21.500 19.000 ;
        RECT 11.500 18.000 22.000 18.500 ;
        RECT 12.000 17.500 22.500 18.000 ;
        RECT 12.500 17.000 23.000 17.500 ;
        RECT 12.500 16.500 24.000 17.000 ;
        RECT 13.000 16.000 24.500 16.500 ;
        RECT 13.500 15.500 25.000 16.000 ;
        RECT 14.000 15.000 26.000 15.500 ;
        RECT 14.500 14.500 26.500 15.000 ;
        RECT 15.000 14.000 27.500 14.500 ;
        RECT 15.500 13.500 28.000 14.000 ;
        RECT 16.000 13.000 29.000 13.500 ;
        RECT 16.500 12.500 30.000 13.000 ;
        RECT 17.500 12.000 31.000 12.500 ;
        RECT 18.000 11.500 32.000 12.000 ;
        RECT 18.500 11.000 33.000 11.500 ;
        RECT 19.000 10.500 34.000 11.000 ;
        RECT 19.500 10.000 35.500 10.500 ;
        RECT 20.500 9.500 37.000 10.000 ;
        RECT 21.000 9.000 38.500 9.500 ;
        RECT 22.000 8.500 40.500 9.000 ;
        RECT 22.500 8.000 43.000 8.500 ;
        RECT 53.500 8.000 68.000 40.500 ;
        RECT 91.000 39.000 99.000 40.500 ;
        RECT 91.000 38.500 98.500 39.000 ;
        RECT 90.500 37.000 98.500 38.500 ;
        RECT 90.000 35.500 98.000 37.000 ;
        RECT 89.500 35.000 98.000 35.500 ;
        RECT 89.500 34.000 97.500 35.000 ;
        RECT 89.000 33.500 97.500 34.000 ;
        RECT 89.000 33.000 97.000 33.500 ;
        RECT 88.500 32.500 97.000 33.000 ;
        RECT 88.500 32.000 96.500 32.500 ;
        RECT 88.000 31.000 96.500 32.000 ;
        RECT 87.500 30.000 96.000 31.000 ;
        RECT 87.000 29.000 95.500 30.000 ;
        RECT 86.500 28.000 95.000 29.000 ;
        RECT 86.000 27.500 94.500 28.000 ;
        RECT 85.500 26.500 94.500 27.500 ;
        RECT 85.000 26.000 94.000 26.500 ;
        RECT 84.500 25.000 93.500 26.000 ;
        RECT 84.000 24.500 93.000 25.000 ;
        RECT 83.500 24.000 93.000 24.500 ;
        RECT 83.000 23.500 92.500 24.000 ;
        RECT 83.000 23.000 92.000 23.500 ;
        RECT 82.500 22.500 92.000 23.000 ;
        RECT 82.000 22.000 91.500 22.500 ;
        RECT 81.500 21.500 91.000 22.000 ;
        RECT 81.000 21.000 91.000 21.500 ;
        RECT 80.500 20.500 90.500 21.000 ;
        RECT 80.000 20.000 90.000 20.500 ;
        RECT 79.500 19.500 90.000 20.000 ;
        RECT 79.000 19.000 89.500 19.500 ;
        RECT 78.500 18.500 89.000 19.000 ;
        RECT 78.000 18.000 88.500 18.500 ;
        RECT 77.500 17.500 88.000 18.000 ;
        RECT 77.000 17.000 87.500 17.500 ;
        RECT 76.000 16.500 87.500 17.000 ;
        RECT 75.500 16.000 87.000 16.500 ;
        RECT 75.000 15.500 86.500 16.000 ;
        RECT 74.000 15.000 86.000 15.500 ;
        RECT 73.500 14.500 85.500 15.000 ;
        RECT 73.000 14.000 85.000 14.500 ;
        RECT 23.500 7.500 47.000 8.000 ;
        RECT 53.000 7.500 68.000 8.000 ;
        RECT 24.000 7.000 68.000 7.500 ;
        RECT 25.000 6.500 68.000 7.000 ;
        RECT 72.500 13.500 84.500 14.000 ;
        RECT 72.500 13.000 84.000 13.500 ;
        RECT 72.500 12.500 83.500 13.000 ;
        RECT 72.500 12.000 83.000 12.500 ;
        RECT 72.500 11.500 82.000 12.000 ;
        RECT 72.500 11.000 81.500 11.500 ;
        RECT 72.500 10.500 81.000 11.000 ;
        RECT 72.500 10.000 80.500 10.500 ;
        RECT 72.500 9.500 79.500 10.000 ;
        RECT 72.500 9.000 79.000 9.500 ;
        RECT 72.500 8.500 78.500 9.000 ;
        RECT 72.500 8.000 77.500 8.500 ;
        RECT 72.500 7.500 76.500 8.000 ;
        RECT 72.500 7.000 76.000 7.500 ;
        RECT 72.500 6.500 75.000 7.000 ;
        RECT 26.000 6.000 68.000 6.500 ;
        RECT 27.000 5.500 68.000 6.000 ;
        RECT 27.500 5.000 68.000 5.500 ;
        RECT 28.500 4.500 68.000 5.000 ;
        RECT 30.000 4.000 68.000 4.500 ;
        RECT 31.000 3.500 68.000 4.000 ;
        RECT 32.500 3.000 67.500 3.500 ;
        RECT 33.500 2.500 66.500 3.000 ;
        RECT 35.000 2.000 65.000 2.500 ;
        RECT 37.000 1.500 63.000 2.000 ;
        RECT 39.000 1.000 61.000 1.500 ;
        RECT 41.500 0.500 58.500 1.000 ;
        RECT 45.000 0.000 55.000 0.500 ;
  END
END tt_logo_corner
END LIBRARY

