`default_nettype none

module tt_logo_top ();
endmodule
